library IEEE;
use IEEE.std_logic_1164.all;

-- Read-phase controller (AR -> R).
-- FSM matches the diagram:
--   s_idle: wait for i_start
--   s_ar  : assert ARVALID until ARREADY handshake
--   s_r   : assert RREADY; finish when last R beat (RVALID&RREADY&RLAST)
--
-- Pulses:
--  * o_txn_start_pulse : 1 cycle when a new transaction starts (IDLE->AR) (registered)
--  * o_rbeat_pulse     : combinational, asserted when R beat is accepted (RVALID&RREADY)
--  * o_done            : 1 cycle when last R beat is accepted (registered)
entity tm_read_controller is
  port(
    ACLK    : in  std_logic;
    ARESETn : in  std_logic := '1';

    -- sequencing
    i_start : in  std_logic := '1';  -- pulse or level; if held '1' it will restart immediately after done
    o_done  : out std_logic;

    -- Handshake inputs (from AXI slave)
    ARREADY : in  std_logic;
    RVALID  : in  std_logic;
    RLAST   : in  std_logic;

    -- AXI control outputs (to AXI slave)
    ARVALID : out std_logic;
    RREADY  : out std_logic;

    -- datapath control
    o_txn_start_pulse : out std_logic;
    o_rbeat_pulse     : out std_logic
  );
end entity;

architecture rtl of tm_read_controller is
  type t_state is (s_idle, s_ar, s_r);
  signal r_state : t_state := s_idle;

  signal arvalid_i, rready_i : std_logic;
  signal ar_hs, r_hs         : std_logic;

  signal done_pulse  : std_logic := '0';
  signal start_pulse : std_logic := '0';
begin
  -- outputs by state
  arvalid_i <= '1' when (r_state = s_ar) else '0';
  rready_i  <= '1' when (r_state = s_r)  else '0';

  ARVALID <= arvalid_i;
  RREADY  <= rready_i;

  -- handshakes
  ar_hs <= arvalid_i and ARREADY;
  r_hs  <= rready_i  and RVALID;

  -- pulses
  o_done            <= done_pulse;
  o_txn_start_pulse <= start_pulse;

  -- IMPORTANT FIX:
  -- rbeat pulse must be asserted in the SAME cycle as the accepted beat,
  -- otherwise the comparator sees RDATA too late.
  o_rbeat_pulse     <= r_hs;

  process(ACLK)
  begin
    if rising_edge(ACLK) then
      done_pulse  <= '0';
      start_pulse <= '0';

      if ARESETn = '0' then
        r_state <= s_idle;
      else
        case r_state is
          when s_idle =>
            if i_start = '1' then
              start_pulse <= '1';
              r_state <= s_ar;
            end if;

          when s_ar =>
            if ar_hs = '1' then
              r_state <= s_r;
            end if;

          when s_r =>
            if r_hs = '1' then
              if RLAST = '1' then
                done_pulse <= '1';
                r_state <= s_idle;
              end if;
            end if;

        end case;
      end if;
    end if;
  end process;

end rtl;
