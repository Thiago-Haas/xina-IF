library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.xina_ft_pkg.all;
use work.xina_ni_ft_pkg.all;

-- TB: TG write manager -> NI manager, with a simple NoC-side loopback.
--
-- Key points (matches the *working* TB behaviour you posted):
--  * lin_ack is a 1-cycle PULSE per accepted flit (this interface behaves like VALID/ACK).
--  * request packet is captured until a flit with ctrl='1' is seen (checksum delimiter).
--  * response is generated by swapping hdr0/hdr1 and rebuilding hdr2.
--
-- Response shaping (aligned with manager_loopback_datapath/tx_response_ctrl):
--  * WRITE response: hdr0, hdr1, hdr2, checksum (NO payload), checksum word = 0x00000000
--  * READ  response: hdr0, hdr1, hdr2, payload[0..LEN], checksum (not used in this TG-write TB)

entity tb_tg_ni_manager_loopback_dbg is
end entity;

architecture tb of tb_tg_ni_manager_loopback_dbg is

  constant c_CLK_PERIOD : time := 10 ns;

  -- multi-transaction regression
  constant c_NUM_ITERS      : natural := 20;
  constant c_TIMEOUT_CYCLES : natural := 50000;

  signal ACLK    : std_logic := '0';
  signal ARESETn : std_logic := '0';

  -- TG control
  signal tg_start : std_logic := '0';
  signal tg_done  : std_logic;
  signal input_address : std_logic_vector(63 downto 0) := (others => '0');
  signal starting_seed : std_logic_vector(31 downto 0) := (others => '0');

  -- NoC side (NI injection = lin_*, NI ejection = lout_*)
  signal lin_data : std_logic_vector(c_FLIT_WIDTH - 1 downto 0);
  signal lin_val  : std_logic;
  signal lin_ack  : std_logic := '0';  -- IMPORTANT: pulse per flit

  signal lout_data : std_logic_vector(c_FLIT_WIDTH - 1 downto 0) := (others => '0');
  signal lout_val  : std_logic := '0';
  signal lout_ack  : std_logic;

  -- ------------------------------------------------------------------
  -- Debug signals exported by tg_ni_write_only_top_dbg
  -- ------------------------------------------------------------------
  signal dbg_axi_awid    : std_logic_vector(c_AXI_ID_WIDTH - 1 downto 0);
  signal dbg_axi_awaddr  : std_logic_vector(c_AXI_ADDR_WIDTH - 1 downto 0);
  signal dbg_axi_awlen   : std_logic_vector(7 downto 0);
  signal dbg_axi_awburst : std_logic_vector(1 downto 0);
  signal dbg_axi_awvalid : std_logic;
  signal dbg_axi_awready : std_logic;

  signal dbg_axi_wvalid  : std_logic;
  signal dbg_axi_wready  : std_logic;
  signal dbg_axi_wdata   : std_logic_vector(c_AXI_DATA_WIDTH - 1 downto 0);
  signal dbg_axi_wlast   : std_logic;

  signal dbg_axi_bid     : std_logic_vector(c_AXI_ID_WIDTH - 1 downto 0);
  signal dbg_axi_bresp   : std_logic_vector(c_AXI_RESP_WIDTH - 1 downto 0);
  signal dbg_axi_bvalid  : std_logic;
  signal dbg_axi_bready  : std_logic;

  signal dbg_tg_state        : std_logic_vector(1 downto 0);
  signal dbg_tg_aw_hs        : std_logic;
  signal dbg_tg_w_hs         : std_logic;
  signal dbg_tg_b_hs         : std_logic;
  signal dbg_tg_bhs_seen     : std_logic;
  signal dbg_tg_txn_start_pulse : std_logic;
  signal dbg_tg_wbeat_pulse     : std_logic;

  signal dbg_dp_seeded       : std_logic;
  signal dbg_dp_do_init      : std_logic;
  signal dbg_dp_do_step      : std_logic;
  signal dbg_dp_init_value   : std_logic_vector(c_AXI_DATA_WIDTH - 1 downto 0);
  signal dbg_dp_feedback_val : std_logic_vector(c_AXI_DATA_WIDTH - 1 downto 0);
  signal dbg_dp_lfsr_input   : std_logic_vector(c_AXI_DATA_WIDTH - 1 downto 0);
  signal dbg_dp_lfsr_next    : std_logic_vector(c_AXI_DATA_WIDTH - 1 downto 0);
  signal dbg_dp_lfsr_in_reg  : std_logic_vector(c_AXI_DATA_WIDTH - 1 downto 0);
  signal dbg_dp_wdata_reg    : std_logic_vector(c_AXI_DATA_WIDTH - 1 downto 0);

  signal dbg_tg_lfsr_value   : std_logic_vector(c_AXI_DATA_WIDTH - 1 downto 0);

  signal dbg_corrupt_packet  : std_logic;

  -- hdr2 bit positions (match manager_loopback_datapath defaults)
  constant c_TYPE_BIT   : integer := 0;
  constant c_OP_BIT     : integer := 1;
  constant c_STATUS_LSB : integer := 2;
  constant c_STATUS_MSB : integer := 3;
  constant c_LENGTH_LSB : integer := 6;
  constant c_LENGTH_MSB : integer := 13;

  -- flit helpers
  function mk_flit(ctrl : std_logic; w : std_logic_vector(31 downto 0)) return std_logic_vector is
    variable f : std_logic_vector(c_FLIT_WIDTH - 1 downto 0) := (others => '0');
  begin
    f(f'left) := ctrl;           -- ctrl at MSB
    f(31 downto 0) := w;
    return f;
  end function;

  subtype t_flit is std_logic_vector(c_FLIT_WIDTH - 1 downto 0);
  constant c_MAX_FLITS : natural := 16; -- enough for small payload tests
  type t_pkt is array(0 to c_MAX_FLITS-1) of t_flit;

  function flit_ctrl(f : t_flit) return std_logic is
  begin
    return f(f'left);
  end function;

  
---------------------------------------------------------------------------
-- Diagnostics helpers
---------------------------------------------------------------------------
constant c_DIAG_ENABLE : boolean := true;
constant c_DIAG_DUMP_PKTS : boolean := true; -- dump every captured packet flit-by-flit

-- 32-bit hex formatting (no std_logic_textio dependency)
function hex32(v : std_logic_vector(31 downto 0)) return string is
  constant H : string := "0123456789ABCDEF";
  variable r : string(1 to 8);
  variable nib : unsigned(3 downto 0);
begin
  for i in 0 to 7 loop
    nib := unsigned(v(31 - i*4 downto 28 - i*4));
    r(i+1) := H(to_integer(nib) + 1);
  end loop;
  return r;
end function;

  -- Format arbitrary std_logic_vector as hex by printing the lower 32 bits (and upper 32 if present).
  function hex_lo32(v : std_logic_vector) return string is
    variable lo : std_logic_vector(31 downto 0) := (others => '0');
  begin
    if v'length >= 32 then
      lo := v(31 downto 0);
    else
      lo(v'length-1 downto 0) := v;
    end if;
    return hex32(lo);
  end function;

  function hex_hi32(v : std_logic_vector) return string is
    variable hi : std_logic_vector(31 downto 0) := (others => '0');
  begin
    if v'length > 32 then
      hi := v(v'length-1 downto 32);
    end if;
    return hex32(hi);
  end function;

procedure dbg(constant msg : in string) is
begin
  if c_DIAG_ENABLE then
    report "t=" & time'image(now) & "  " & msg severity note;
  end if;
end procedure;

procedure dump_flit(constant tag : in string; constant idx : in natural; constant f : in t_flit) is
begin
  if c_DIAG_ENABLE then
    report "t=" & time'image(now) & "  " & tag &
           " [" & integer'image(integer(idx)) & "] ctrl=" & std_logic'image(f(f'left)) &
           " word=0x" & hex32(f(31 downto 0))
      severity note;
  end if;
end procedure;

function set_bit(v : std_logic_vector(31 downto 0); idx : integer; b : std_logic) return std_logic_vector is
    variable r : std_logic_vector(31 downto 0) := v;
  begin
    r(idx) := b;
    return r;
  end function;

  function set_slice(v : std_logic_vector(31 downto 0); lsb : integer; msb : integer; s : std_logic_vector) return std_logic_vector is
    variable r : std_logic_vector(31 downto 0) := v;
  begin
    r(msb downto lsb) := s;
    return r;
  end function;

  signal sim_done : std_logic := '0';

begin

  -- clock
  ACLK <= not ACLK after c_CLK_PERIOD/2;

  -- DUT
  u_dut: entity work.tg_ni_write_only_top_dbg
    port map(
      ACLK    => ACLK,
      ARESETn => ARESETn,

      i_start       => tg_start,
      o_done        => tg_done,
      INPUT_ADDRESS => input_address,
      STARTING_SEED => starting_seed,

      l_in_data_o => lin_data,
      l_in_val_o  => lin_val,
      l_in_ack_i  => lin_ack,

      l_out_data_i => lout_data,
      l_out_val_i  => lout_val,
      l_out_ack_o  => lout_ack,

      -- Debug exports
      o_dbg_axi_awid    => dbg_axi_awid,
      o_dbg_axi_awaddr  => dbg_axi_awaddr,
      o_dbg_axi_awlen   => dbg_axi_awlen,
      o_dbg_axi_awburst => dbg_axi_awburst,
      o_dbg_axi_awvalid => dbg_axi_awvalid,
      o_dbg_axi_awready => dbg_axi_awready,

      o_dbg_axi_wvalid  => dbg_axi_wvalid,
      o_dbg_axi_wready  => dbg_axi_wready,
      o_dbg_axi_wdata   => dbg_axi_wdata,
      o_dbg_axi_wlast   => dbg_axi_wlast,

      o_dbg_axi_bid     => dbg_axi_bid,
      o_dbg_axi_bresp   => dbg_axi_bresp,
      o_dbg_axi_bvalid  => dbg_axi_bvalid,
      o_dbg_axi_bready  => dbg_axi_bready,

      o_dbg_tg_state        => dbg_tg_state,
      o_dbg_tg_aw_hs        => dbg_tg_aw_hs,
      o_dbg_tg_w_hs         => dbg_tg_w_hs,
      o_dbg_tg_b_hs         => dbg_tg_b_hs,
      o_dbg_tg_bhs_seen     => dbg_tg_bhs_seen,
      o_dbg_tg_txn_start_pulse => dbg_tg_txn_start_pulse,
      o_dbg_tg_wbeat_pulse     => dbg_tg_wbeat_pulse,

      o_dbg_dp_seeded       => dbg_dp_seeded,
      o_dbg_dp_do_init      => dbg_dp_do_init,
      o_dbg_dp_do_step      => dbg_dp_do_step,
      o_dbg_dp_init_value   => dbg_dp_init_value,
      o_dbg_dp_feedback_val => dbg_dp_feedback_val,
      o_dbg_dp_lfsr_input   => dbg_dp_lfsr_input,
      o_dbg_dp_lfsr_next    => dbg_dp_lfsr_next,
      o_dbg_dp_lfsr_in_reg  => dbg_dp_lfsr_in_reg,
      o_dbg_dp_wdata_reg    => dbg_dp_wdata_reg,

      o_dbg_tg_lfsr_value   => dbg_tg_lfsr_value,

      o_dbg_corrupt_packet  => dbg_corrupt_packet
    );


  ---------------------------------------------------------------------------
  -- AXI/TG/NI monitor (prints state changes, handshakes, and a periodic snapshot)
  ---------------------------------------------------------------------------
  monitor: process
    variable prev_state : std_logic_vector(1 downto 0) := (others => 'X');
    variable stall_cnt  : natural := 0;
  begin
    wait until ARESETn = '1';
    wait until rising_edge(ACLK);

    while sim_done = '0' loop
      wait until rising_edge(ACLK);

      -- State transitions
      if dbg_tg_state /= prev_state then
        dbg("TG STATE " & std_logic'image(prev_state(1)) & std_logic'image(prev_state(0)) &
            " -> " & std_logic'image(dbg_tg_state(1)) & std_logic'image(dbg_tg_state(0)) &
            " | AWV/AWR=" & std_logic'image(dbg_axi_awvalid) & "/" & std_logic'image(dbg_axi_awready) &
            " WV/WR=" & std_logic'image(dbg_axi_wvalid) & "/" & std_logic'image(dbg_axi_wready) &
            " BV/BR=" & std_logic'image(dbg_axi_bvalid) & "/" & std_logic'image(dbg_axi_bready) &
            " corrupt=" & std_logic'image(dbg_corrupt_packet));
        prev_state := dbg_tg_state;
      end if;

      -- Handshake event prints (AW/W/B)
      if dbg_tg_aw_hs = '1' then
        dbg("AXI AW_HS: awid=" & integer'image(to_integer(unsigned(dbg_axi_awid))) &
            " awaddr_hi=0x" & hex_hi32(dbg_axi_awaddr) &
            " awaddr_lo=0x" & hex_lo32(dbg_axi_awaddr) &
            " awlen=" & integer'image(to_integer(unsigned(dbg_axi_awlen))) &
            " awburst=" & integer'image(to_integer(unsigned(dbg_axi_awburst))));
      end if;

      if dbg_tg_w_hs = '1' then
        dbg("AXI W_HS: wlast=" & std_logic'image(dbg_axi_wlast) &
            " wdata_hi=0x" & hex_hi32(dbg_axi_wdata) &
            " wdata_lo=0x" & hex_lo32(dbg_axi_wdata) &
            " | seeded=" & std_logic'image(dbg_dp_seeded) &
            " do_init/do_step=" & std_logic'image(dbg_dp_do_init) & "/" & std_logic'image(dbg_dp_do_step) &
            " lfsr_in_lo=0x" & hex_lo32(dbg_dp_lfsr_input) &
            " lfsr_next_lo=0x" & hex_lo32(dbg_dp_lfsr_next));
      end if;

      if dbg_tg_b_hs = '1' then
        dbg("AXI B_HS: bid=" & integer'image(to_integer(unsigned(dbg_axi_bid))) &
            " bresp=" & integer'image(to_integer(unsigned(dbg_axi_bresp))) &
            " bhs_seen=" & std_logic'image(dbg_tg_bhs_seen) &
            " corrupt=" & std_logic'image(dbg_corrupt_packet));
      end if;

      -- Detect NoC activity
      if lin_val = '1' then
        stall_cnt := 0;
      elsif lout_val = '1' then
        stall_cnt := 0;
      else
        stall_cnt := stall_cnt + 1;
      end if;

      if stall_cnt = 2000 then
        dbg("---- STALL SNAPSHOT ----");
        dbg("TG state=" & std_logic'image(dbg_tg_state(1)) & std_logic'image(dbg_tg_state(0)) &
            " AWV/AWR=" & std_logic'image(dbg_axi_awvalid) & "/" & std_logic'image(dbg_axi_awready) &
            " WV/WR=" & std_logic'image(dbg_axi_wvalid) & "/" & std_logic'image(dbg_axi_wready) &
            " BV/BR=" & std_logic'image(dbg_axi_bvalid) & "/" & std_logic'image(dbg_axi_bready));
        dbg("AW: id=" & integer'image(to_integer(unsigned(dbg_axi_awid))) &
            " addr_hi=0x" & hex_hi32(dbg_axi_awaddr) & " addr_lo=0x" & hex_lo32(dbg_axi_awaddr) &
            " len=" & integer'image(to_integer(unsigned(dbg_axi_awlen))) &
            " burst=" & integer'image(to_integer(unsigned(dbg_axi_awburst))));
        dbg("W : last=" & std_logic'image(dbg_axi_wlast) &
            " data_hi=0x" & hex_hi32(dbg_axi_wdata) & " data_lo=0x" & hex_lo32(dbg_axi_wdata));
        dbg("B : valid=" & std_logic'image(dbg_axi_bvalid) &
            " resp=" & integer'image(to_integer(unsigned(dbg_axi_bresp))) &
            " id=" & integer'image(to_integer(unsigned(dbg_axi_bid))));
        dbg("NoC: lin_val=" & std_logic'image(lin_val) & " lin_ack=" & std_logic'image(lin_ack) &
            " | lout_val=" & std_logic'image(lout_val) & " lout_ack=" & std_logic'image(lout_ack));
        dbg("DP : seeded=" & std_logic'image(dbg_dp_seeded) &
            " lfsr_in_reg_lo=0x" & hex_lo32(dbg_dp_lfsr_in_reg) &
            " wdata_reg_lo=0x" & hex_lo32(dbg_dp_wdata_reg));
      end if;
    end loop;
    wait;
  end process;

  ---------------------------------------------------------------------------
  -- NoC loopback emulator
  ---------------------------------------------------------------------------
  noc_loopback: process
    variable req  : t_pkt;
    variable req_len  : natural;

    variable req_hdr0 : std_logic_vector(31 downto 0);
    variable req_hdr1 : std_logic_vector(31 downto 0);
    variable req_hdr2 : std_logic_vector(31 downto 0);

    variable req_type : std_logic;
    variable req_op   : std_logic;
    variable req_len_field : unsigned(7 downto 0);

    variable resp_hdr0 : std_logic_vector(31 downto 0);
    variable resp_hdr1 : std_logic_vector(31 downto 0);
    variable resp_hdr2 : std_logic_vector(31 downto 0);

    variable payload_words : natural;
    variable req_payload_words : natural;

    variable resp_idx : natural;
    variable plw : std_logic_vector(31 downto 0);

    variable cyc : natural;

    -- Accept exactly one outgoing flit (NI->TB): sample, then pulse lin_ack
    -- Accept exactly one outgoing flit (NI->TB): sample, then pulse lin_ack
-- This TB uses the "VALID/ACK pulse" semantics the user described.
procedure accept_one_req_flit(variable dst : out t_flit; constant idx : in natural) is
begin
  cyc := 0;

  -- wait for a flit to appear
  while lin_val /= '1' loop
    wait until rising_edge(ACLK);
    if sim_done = '1' then
      dst := (others => '0');
      return;
    end if;
    cyc := cyc + 1;
    if (cyc mod 1000) = 0 then
      dbg("...waiting lin_val for request flit idx=" & integer'image(integer(idx)) &
          " (cycles waited=" & integer'image(integer(cyc)) & ")");
    end if;
    if cyc = c_TIMEOUT_CYCLES then
      assert false report "TIMEOUT waiting lin_val (request flit)" severity failure;
    end if;
  end loop;

  -- sample with ACK low (NI must hold stable until ACK pulses)
  wait for 1 ns;
  dst := lin_data;
  dump_flit("RX", idx, dst);

  -- pulse ACK for one cycle to advance to next flit
  dbg("PULSE lin_ack for RX idx=" & integer'image(integer(idx)));
  lin_ack <= '1';
  wait until rising_edge(ACLK);
  lin_ack <= '0';
  wait until rising_edge(ACLK);
end procedure;

    -- Send one response flit (TB->NI): hold until NI asserts lout_ack
    -- Send one response flit (TB->NI): hold VAL high until NI asserts lout_ack
procedure send_resp_flit(constant f : in t_flit; constant idx : in natural) is
begin
  dump_flit("TX", idx, f);
  lout_val  <= '1';
  lout_data <= f;
  cyc := 0;
  loop
    wait until rising_edge(ACLK);
    exit when lout_ack = '1';
    cyc := cyc + 1;
    if (cyc mod 1000) = 0 then
      dbg("...waiting lout_ack for response flit idx=" & integer'image(integer(idx)) &
          " (cycles waited=" & integer'image(integer(cyc)) & ")");
    end if;
    if cyc = c_TIMEOUT_CYCLES then
      assert false report "TIMEOUT waiting lout_ack (sending response flit)" severity failure;
    end if;
  end loop;
  dbg("Got lout_ack for TX idx=" & integer'image(integer(idx)));
end procedure;

  begin
    -- init outputs
    lin_ack   <= '0';
    lout_val  <= '0';
    lout_data <= (others => '0');

    wait until ARESETn = '1';
    wait until rising_edge(ACLK);

    while sim_done = '0' loop
      ---------------------------------------------------------------------
      -- Capture one full request packet, stopping on checksum flit (ctrl='1').
      ---------------------------------------------------------------------
      req_len := 0;

      -- hdr0
      accept_one_req_flit(req(0), 0);
      if sim_done = '1' then
        exit;
      end if;
      assert flit_ctrl(req(0)) = '1'
        report "Expected ctrl=1 on hdr0" severity failure;
      req_len := 1;

      -- capture until checksum (ctrl='1')
      while req_len < c_MAX_FLITS loop
        accept_one_req_flit(req(req_len), req_len);
        if sim_done = '1' then
          exit;
        end if;
        req_len := req_len + 1;
        exit when flit_ctrl(req(req_len-1)) = '1';
      end loop;

      assert req_len < c_MAX_FLITS
        report "Request packet too long (no checksum delimiter)" severity failure;


if c_DIAG_DUMP_PKTS then
  dbg("---- BEGIN REQUEST PACKET DUMP (flits=" & integer'image(integer(req_len)) & ") ----");
  for k in 0 to integer(req_len)-1 loop
    dump_flit("REQ", natural(k), req(k));
  end loop;
  dbg("---- END   REQUEST PACKET DUMP ----");

-- Infer whether the REQUEST carries payload (WRITE request has payload flits, READ request doesn't)
-- Minimal request flits = 5 (hdr0,hdr1,hdr2,addr,checksum). Any extra before checksum are payload.
req_payload_words := 0;
if req_len > 5 then
  req_payload_words := req_len - 5;
end if;
dbg("REQ inferred payload_words=" & integer'image(integer(req_payload_words)));

end if;

      -- basic decode (need at least hdr0,hdr1,hdr2)
      assert req_len >= 3
        report "Request packet too short" severity failure;

      req_hdr0 := req(0)(31 downto 0);
      req_hdr1 := req(1)(31 downto 0);
      req_hdr2 := req(2)(31 downto 0);

      req_type := req_hdr2(c_TYPE_BIT);
      req_op   := req_hdr2(c_OP_BIT);
      req_len_field := unsigned(req_hdr2(c_LENGTH_MSB downto c_LENGTH_LSB));

      -- optional info
            report "RX pkt: flits=" & integer'image(integer(req_len)) &
             "  hdr0=0x" & hex32(req_hdr0) &
             "  hdr1=0x" & hex32(req_hdr1) &
             "  hdr2=0x" & hex32(req_hdr2) &
             "  TYPE=" & std_logic'image(req_type) &
             "  OP=" & std_logic'image(req_op) &
             "  LEN=" & integer'image(to_integer(req_len_field))
        severity note;

      ---------------------------------------------------------------------
      -- Build response (swap hdr0/hdr1, force TYPE=1, STATUS=00)
      ---------------------------------------------------------------------
      resp_hdr0 := req_hdr0;
      resp_hdr1 := req_hdr1;

      dbg("RESP build: hdr0=0x" & hex32(resp_hdr0) &
          " hdr1=0x" & hex32(resp_hdr1));

      resp_hdr2 := req_hdr2;
resp_hdr2 := set_bit(resp_hdr2, c_TYPE_BIT, '1');
resp_hdr2 := set_slice(resp_hdr2, c_STATUS_LSB, c_STATUS_MSB, "00");

-- Decide response payload length WITHOUT trusting OP bit positions:
-- If the request carried payload flits => it's a WRITE request => WRITE response has NO payload.
-- Otherwise => it's a READ request => READ response has LEN+1 payload words.
if (req_type = '0') then
  if req_payload_words > 0 then
    -- WRITE response
    payload_words := 0;
    resp_hdr2 := set_slice(resp_hdr2, c_LENGTH_LSB, c_LENGTH_MSB,
                         std_logic_vector(to_unsigned(0, c_LENGTH_MSB-c_LENGTH_LSB+1)));
  else
    -- READ response
    payload_words := to_integer(req_len_field) + 1;
  end if;
else
  -- If it's not a request, default to no payload
  payload_words := 0;
end if;

      ---------------------------------------------------------------------
      -- Send response packet
      --  hdr0(ctrl=1), hdr1, hdr2, [payload], checksum(ctrl=1)
      --  checksum word is ZERO (as in manager_loopback_datapath)
      ---------------------------------------------------------------------
      resp_idx := 0;

-- Response format must match tx_response_ctrl:
--   hdr0, hdr1, hdr2, [payload words if READ], checksum
--   (No address flit is transmitted in the response.)
--
-- hdr0
send_resp_flit(mk_flit('1', resp_hdr0), resp_idx);
resp_idx := resp_idx + 1;

-- hdr1
send_resp_flit(mk_flit('0', resp_hdr1), resp_idx);
resp_idx := resp_idx + 1;

-- hdr2
send_resp_flit(mk_flit('0', resp_hdr2), resp_idx);
resp_idx := resp_idx + 1;

-- payload (only when payload_words > 0): send that many words
if payload_words > 0 then
  -- We don't have real memory here; return a deterministic word so the NI can complete.
  -- If there was at least one extra captured flit after addr, echo it; else return 0.
  plw := (others => '0');
  if req_len > 5 then
    plw := req(4)(31 downto 0);
  end if;

  for p in 0 to integer(payload_words)-1 loop
    send_resp_flit(mk_flit('0', plw), resp_idx);
    resp_idx := resp_idx + 1;
  end loop;
end if;

-- checksum
send_resp_flit(mk_flit('1', (others => '0')), resp_idx);
resp_idx := resp_idx + 1;

      -- release bus
      lout_val  <= '0';
      lout_data <= (others => '0');
      wait until rising_edge(ACLK);

    end loop;

    -- clean
    lout_val  <= '0';
    lout_data <= (others => '0');
    lin_ack   <= '0';
    wait;
  end process;

  ---------------------------------------------------------------------------
  -- Stimulus: multiple GO iterations
  ---------------------------------------------------------------------------
  stim: process
    variable cyc : natural;
  begin
    tg_start      <= '0';
    input_address <= x"0000_0000_0000_0100";
    starting_seed <= x"1ACE_B00C";

    -- reset
    ARESETn <= '0';
    wait for 100 ns;
    wait until rising_edge(ACLK);
    ARESETn <= '1';
    wait until rising_edge(ACLK);

    for it in 0 to integer(c_NUM_ITERS)-1 loop
      dbg("=== ITER " & integer'image(it) & " START: addr=0x" & hex32(input_address(31 downto 0)) & " seed=0x" & hex32(starting_seed) & " ===");
      -- pulse start (1 cycle)
      tg_start <= '1';
      wait until rising_edge(ACLK);
      tg_start <= '0';

      -- wait done
      cyc := 0;
      while tg_done /= '1' loop
        wait until rising_edge(ACLK);
        cyc := cyc + 1;
        if cyc = c_TIMEOUT_CYCLES then
          assert false report "TIMEOUT waiting tg_done at iter=" & integer'image(it) severity failure;
        end if;
      end loop;

      dbg("=== ITER " & integer'image(it) & " DONE (tg_done seen) ===");
      -- small gap
      wait until rising_edge(ACLK);
      wait until rising_edge(ACLK);

      -- vary address/seed
      input_address <= std_logic_vector(unsigned(input_address) + 16);
      starting_seed <= std_logic_vector(unsigned(starting_seed) + 1);
    end loop;

    sim_done <= '1';
    report "TB completed OK" severity note;
    wait for 50 ns;
    assert false report "End of simulation" severity failure;
  end process;

end architecture;
